`include "uvm_macros.svh"
import uvm_pkg::*;

class cic_filter_transaction extends uvm_sequence_item;
  `uvm_object_utils(cic_filter_transaction)

  bit [15:0] data;

  // Construtor deve ser definido aqui

endclass

