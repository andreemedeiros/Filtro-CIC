`include "uvm_macros.svh"
import uvm_pkg::*;
`include "cic_filter_transaction.sv"

class cic_filter_scoreboard extends uvm_scoreboard;
  `uvm_component_utils(cic_filter_scoreboard)

  // Construtor e outros métodos devem ser definidos aqui

endclass
